library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;


entity ControlFlow is
	generic (
		ADDR_WIDTH : integer := 8;	
		DATA_WIDTH : integer := 32
	);
	port (
		clk, reset : in std_logic;
		pc_out : out std_logic_vector(ADDR_WIDTH-1 downto 0);
		instruction_in : in std_logic_vector(DATA_WIDTH-1 downto 0);
		alu_zero_in, branch_in, jump_in, pc_write_in : in std_logic
	);

end ControlFlow;

architecture Behavioral of ControlFlow is

	signal pc, pc_in, pc_add_1, pc_jump, pc_immediate_signextend, pc_add_immediate, pc_branch : signed(DATA_WIDTH-1 downto 0);
	
begin

	-- Process for PC register
	PCBehaviour: process(clk, reset)
	begin
		if reset = '1' then
			pc <= (others => '0');
		elsif rising_edge(clk) and pc_write_in = '1' then
			-- Handle Jumps
			if jump_in = '1' then
				pc <= (pc and "11111100000000000000000000000000") or (signed(instruction_in) and "00000011111111111111111111111111");
			-- Handle branches
			elsif branch_in = '1' and alu_zero_in = '1' then
				pc <= pc + 1 + resize(signed(instruction_in(15 downto 0)), DATA_WIDTH);
			-- Handle increment by 1
			else
				pc <= pc + 1;
			end if;
		end if;
	end process;
	pc_out <= std_logic_vector(pc(ADDR_WIDTH-1 downto 0));



end Behavioral;

